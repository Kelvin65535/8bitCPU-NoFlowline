library ieee;
use ieee.std_logic_1164.all;

---------------AR��ַ�Ĵ���---------------
--���Ҫ��д���ڴ浥Ԫ�ĵ�ַ

--��Ҫִ��ָ��ʱ��ָ��ĵ�ַ��ӳ��������ת��AR��ַ�Ĵ���Ȼ��PC����1
--����û��cache�����PC��ֱ�Ӵ�ŵ�ַ����ֱ���͵�AR
--��AR��ַ�Ĵ����ѵ�ַ���͵���ַ����
--��ַ���߻���յ�ַ���ѵ�ַ��Ӧ���ڴ浥Ԫ������ͨ���������߷��͵�IRָ��Ĵ���

--�������Ϊ����PC��������������ĵ�ַ������ALU������Զ�д�ڴ�ָ��ĵ�ַ
--���Ϊ��Ҫ���ʵĵ�ַ�������Ǵ��ڴ浥Ԫ��ȡ��������ݣ���������ַ����

--��IR��ָ��Ĵ��������ÿ����ź�REC

--------------REC�����ź�˵��--------------
------|REC|--------|      ����      |-----
------|---|--------|----------------|-----
------| 00|--------|     �޲���     |-----
------| 01|--------| AR����PC�ĵ�ַ  |-----
------| 11|--------| AR����ALU����� |-----
------| 10|--------|   AR��������    |-----
------------------------------------------

----ʵ��˵��----
entity ar is
	port(
		 --��alu_out���վ���ALU�����ĵ�ַ
		 alu_out:   in std_logic_vector(7 downto 0);
	     --��pc��������pc����������ĵ�ַ
	     pc:        in std_logic_vector(7 downto 0);
	     --recΪAR����������Դ�Ŀ����ź�
	     rec:       in std_logic_vector(1 downto 0);
	     --clkΪʱ�ӣ�resetΪ��λ��reset�͵�ƽ��Ч
	     clk,reset: in std_logic;
	     --qΪ�����ַ��������ַ����
	     q:         out std_logic_vector(15 downto 0));
end ar;

----ʵ����Ϊ˵��----
architecture behave of ar is
begin
	process(clk,reset)
	begin
		--��resetΪ�͵�ƽʱAR�Ĵ�������
		if reset = '0' then            
        	q <= "0000000000000000";
        --��ʱ������������ʱ����AR����
        elsif clk'event and clk = '1' then
			--ͨ��rec�����ź�ѡ��AR���յ�ַ����Դ
			case rec is
				--��recΪ01ʱ��PC������������յ�ַ
				when "01"=>
					q <= "00000000" & pc;
				--��recΪ11ʱ��ALU���յ�ַ
				when "11"=>
					q <= "00000000" & alu_out;
				--���������ʱAR��������
				when others=>
					null;
			end case;		
        end if;
	end process;
end behave;